// alu testbench
module alu #(
  parameter int W = 4
)
  input
